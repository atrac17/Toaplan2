/*
* <-- pr4m0d -->
* https://pram0d.com
* https://twitter.com/pr4m0d
* https://github.com/psomashekar
*
* Copyright (c) 2022 Pramod Somashekar
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU General Public License as published by
* the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU General Public License for more details.
*
* You should have received a copy of the GNU General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
*/
module snowbro2_game(
    //clock and reset
    input rst,
    input rst48,
    input rst96,
    input rst24, //27mhz
    input rst6, //6.75mhz
    input clk,
    input clk48,
    input clk96,
    input clk24,
    input clk6,
    output pxl_cen,
    output pxl2_cen,

    //video outputs
    output [7:0] red,
    output [7:0] green,
    output [7:0] blue,
    output LHBL,
    output LVBL,
    output HS,
    output VS,

    // Control I/O
    input [3:0] start_button,
    input [3:0] coin_input,
    input [9:0] joystick1,
    input [9:0] joystick2,
    input [9:0] joystick3,
    input [9:0] joystick4,

    // SDRAM interface
    output [21:0] ba0_addr,
    output [21:0] ba1_addr,
    output [21:0] ba2_addr,
    output [21:0] ba3_addr,
    output  [3:0] ba_rd,
    output        ba_wr,
    output [15:0] ba0_din,
    output  [1:0] ba0_din_m,
    input   [3:0] ba_ack,
    input   [3:0] ba_dst,
    input   [3:0] ba_dok,
    input   [3:0] ba_rdy,
    input  [15:0] data_read,

    //ROM loader
    input         downloading,
    output        dwnld_busy,
    input  [25:0] ioctl_addr,
    input   [7:0] ioctl_dout,
    input         ioctl_wr,
    output  [7:0] ioctl_din,
    input         ioctl_ram,
    output [21:0] prog_addr,
    output [15:0] prog_data,
    output  [1:0] prog_mask,
    output  [1:0] prog_ba,
    output        prog_we,
    output        prog_rd,
    input         prog_ack,
    input         prog_dok,
    input         prog_dst,
    input         prog_rdy,

    //dip switches
    input [31:0] status,
    input        service,
    input        dip_pause,
    inout        dip_flip,
    input        dip_test,
    input  [1:0] dip_fxlevel,
    input [31:0] dipsw,

    //sound
    output signed [15:0] snd_left,
    output signed [15:0] snd_right,
    output               sample,
    input                enable_psg,
    input                enable_fm,

    //misc
    output       game_led,
    output       user_led,
    input        gfx_en
);

/*MAIN GLOBALS*/
localparam DEFAULT = 0, SNOWBRO2 = 2;
wire RESET = rst48;
wire CLK = clk48;
wire CLK96 = clk;
wire CLK24 = clk24;
wire CLK6 = clk6;
wire RESET96 = rst;
wire RESET24 = rst24;
wire RESET6 = rst6;

wire CEN16, CEN16B;
wire FLIP = GAME==DEFAULT  ? dipsw[1]:  // Placeholder
            GAME==SNOWBRO2 ? dipsw[1]:  // Screen inversion for SNOWBRO2
            0;

// assign game_led = downloading ? 1'b0 : 1'b1;

/*CLOCKS*/
wire CEN675, CEN675B, CEN2p7, CEN2p7B, CEN1350, CEN1350B;
wire CEN3p375, CEN3p375B, CEN1p6875, CEN1p6875B;
snowbro2_clock u_clocken (
    .CLK(CLK),
    .CLK96(CLK96),
    .CLK24(CLK24),
    .CLK6(CLK6),
    .CEN675(CEN675),
    .CEN675B(CEN675B),
    .CEN2p7(CEN2p7),
    .CEN2p7B(CEN2p7B),
    .CEN3p375(CEN3p375),
    .CEN3p375B(CEN3p375B),
    .CEN1p6875(CEN1p6875),
    .CEN1p6875B(CEN1p6875B),
    .CEN1350(CEN1350),
    .CEN1350B(CEN1350B)
);

assign pxl_cen = CEN675;
assign pxl2_cen = CEN1350;

/*MEMORY CONNECTS*/
//GAME selector
wire [7:0] GAME;
//68K ROM
wire ROM68K_CS;
wire ROM68K_OK;
wire [18:0] ROM68K_ADDR;
wire [15:0] ROM68K_DOUT;

//sound
wire                YM2151_CS;
wire                OKI_CS;
wire                YM2151_WE;
wire                YM2151_WR_CMD;
wire                OKI_WE;
wire          [7:0] OKI_DIN;
wire          [7:0] YM2151_DIN;
wire          [7:0] YM2151_DOUT;
wire          [7:0] OKI_DOUT;
wire                OKI_BANK;
wire                YM2151_INT;

//PCM
wire PCM_CS;
wire PCM_OK;
wire  [19:0] PCM_ADDR;
wire  [7:0]  PCM_DOUT;

//TILE GFX ROM
wire  GFX_CS;
wire  GFX_OK;
wire [21:0] GFX0_ADDR;
wire [31:0] GFX0_DOUT;

wire  GFXSCR0_CS;
wire  GFXSCR0_OK;
wire [21:0] GFX0SCR0_ADDR;
wire [31:0] GFX0SCR0_DOUT;

wire  GFXSCR1_CS;
wire  GFXSCR1_OK;
wire [21:0] GFX0SCR1_ADDR;
wire [31:0] GFX0SCR1_DOUT;

wire  GFXSCR2_CS;
wire  GFXSCR2_OK;
wire [21:0] GFX0SCR2_ADDR;
wire [31:0] GFX0SCR2_DOUT;

//EEPROM
wire EEPROM_SCLK, EEPROM_SCS, EEPROM_SDI, EEPROM_SDO;

/*EXTERNAL DEVICES*/

//gp9001
wire GP9001ACK;
wire GP9001CS, VINT;
wire GP9001_OP_SELECT_REG, GP9001_OP_WRITE_REG, GP9001_OP_WRITE_RAM, GP9001_OP_READ_RAM_H, GP9001_OP_READ_RAM_L, GP9001_OP_SET_RAM_PTR, GP9001_OP_OBJECTBANK_WR;
wire [2:0] GP9001_OBJECTBANK_SLOT;
wire [15:0] CPU_DOUT;
wire [15:0] GCU_DOUT;
wire [10:0] GP9001OUT;

//bus sharing
wire BUSACK;
wire BR = 1'b0;

//dip switch
wire [23:0] DIPSW = GAME == DEFAULT ? {dipsw[23:2], 1'b0, dipsw[0]} :    // Placeholder
                    GAME == SNOWBRO2 ? {dipsw[23:2], 1'b0, dipsw[0]} :   // Screen inversion for SNOWBRO2
                    dipsw[23:0];
wire DIP_TEST = dip_test;
wire DIP_PAUSE = dip_pause;
wire [7:0] DIPSW_C, DIPSW_B, DIPSW_A;
assign { DIPSW_C, DIPSW_B, DIPSW_A } = DIPSW[23:0];

//video timings
wire HSYNC, VSYNC, FBLANK;
wire LHBLL, LVBLL;
wire [8:0] V;

//vrams
wire [10:0] PALRAM_ADDR;
wire [15:0] PALRAM_DATA;
wire [13:0] SRAM_ADDR;
wire [7:0] SRAM_DATA;
wire [7:0] SRAM_DIN;
wire SRAM_WE;


    //cpu
snowbro2_cpu u_cpu (
    .CLK(CLK),
    .CLK96(CLK96),
    .CEN16(CEN16),
    .CEN16B(CEN16B),
    .BUSACK(BUSACK),
    .BR(BR),
    .RESET(RESET),
    .RESET96(RESET96),
    .DOUT(CPU_DOUT),
    .LVBL(LVBLL), //this is low active to the CPU
    .V(V),
    .FLIP(FLIP),

    //inputs
    .JOYMODE(0),
    .JOYSTICK1(joystick1),
    .JOYSTICK2(joystick2),
    .JOYSTICK3(joystick3),
    .JOYSTICK4(joystick4),
    .START_BUTTON(start_button),
    .COIN_INPUT(coin_input),
    .SERVICE(service),
    .TILT(1'b0),

    //dip switches
    .DIPSW_A(DIPSW_A),
    .DIPSW_B(DIPSW_B),
    .DIPSW_C(DIPSW_C),
    .DIP_TEST(DIP_TEST),
    .DIP_PAUSE(DIP_PAUSE),

    //68k program
    .CPU_PRG_CS(ROM68K_CS),
    .CPU_PRG_OK(ROM68K_OK),
    .CPU_PRG_ADDR(ROM68K_ADDR), //16bit addressing
    .CPU_PRG_DATA(ROM68K_DOUT),

    //gcu communications
    .GP9001CS(GP9001CS),
    .GP9001ACK(GP9001ACK),
    .VINT(VINT),
    .GP9001_OP_SELECT_REG(GP9001_OP_SELECT_REG),
    .GP9001_OP_WRITE_REG(GP9001_OP_WRITE_REG),
    .GP9001_OP_WRITE_RAM(GP9001_OP_WRITE_RAM),
    .GP9001_OP_READ_RAM_H(GP9001_OP_READ_RAM_H),
    .GP9001_OP_READ_RAM_L(GP9001_OP_READ_RAM_L),
    .GP9001_OP_SET_RAM_PTR(GP9001_OP_SET_RAM_PTR),
    .GP9001_DOUT(GCU_DOUT),
    .HSYNC(HSYNC),
    .VSYNC(VSYNC),
    .FBLANK(FBLANK),

    //VRAMs
    .PALRAM_ADDR(PALRAM_ADDR),
    .PALRAM_DATA(PALRAM_DATA),

    .GAME(GAME),

    //sound communications
    .YM2151_CS(YM2151_CS),
    .OKI_CS(OKI_CS),
    .YM2151_WE(YM2151_WE),
    .YM2151_WR_CMD(YM2151_WR_CMD),
    .OKI_WE(OKI_WE),
    .OKI_DIN(OKI_DIN),
    .YM2151_DIN(YM2151_DIN),
    .YM2151_DOUT(YM2151_DOUT),
    .OKI_DOUT(OKI_DOUT),
    .OKI_BANK(OKI_BANK),
    .YM2151_INT(YM2151_INT)
);

raizing_video u_video(
    .CLK(CLK),
    .CLK96(CLK96),
    .PIXEL_CEN(pxl_cen),
    .RESET(RESET),
    .RESET96(RESET96),

    //graphics ROM
    .GFX_CS(GFX_CS),
    .GFX_OK(GFX_OK),
    .GFX0_ADDR(GFX0_ADDR),
    .GFX0_DOUT(GFX0_DOUT),

    .GFXSCR0_CS(GFXSCR0_CS),
    .GFXSCR0_OK(GFXSCR0_OK),
    .GFX0SCR0_ADDR(GFX0SCR0_ADDR),
    .GFX0SCR0_DOUT(GFX0SCR0_DOUT),

    .GFXSCR1_CS(GFXSCR1_CS),
    .GFXSCR1_OK(GFXSCR1_OK),
    .GFX0SCR1_ADDR(GFX0SCR1_ADDR),
    .GFX0SCR1_DOUT(GFX0SCR1_DOUT),

    .GFXSCR2_CS(GFXSCR2_CS),
    .GFXSCR2_OK(GFXSCR2_OK),
    .GFX0SCR2_ADDR(GFX0SCR2_ADDR),
    .GFX0SCR2_DOUT(GFX0SCR2_DOUT),

    //gp9001
    .GP9001CS(GP9001CS),
    .GP9001ACK(GP9001ACK),
    .VINT(VINT),
    .GP9001DIN(CPU_DOUT),
    .GP9001DOUT(GCU_DOUT),
    .GP9001_OP_SELECT_REG(GP9001_OP_SELECT_REG),
    .GP9001_OP_WRITE_REG(GP9001_OP_WRITE_REG),
    .GP9001_OP_WRITE_RAM(GP9001_OP_WRITE_RAM),
    .GP9001_OP_READ_RAM_H(GP9001_OP_READ_RAM_H),
    .GP9001_OP_READ_RAM_L(GP9001_OP_READ_RAM_L),
    .GP9001_OP_SET_RAM_PTR(GP9001_OP_SET_RAM_PTR),
    .GP9001OUT(GP9001OUT),

    //video signal
    .LVBL_DLY(LVBL),
    .LHBL_DLY(LHBL),
    .LVBL(LVBLL),
    .LHBL(LHBLL),
    .HS(HS),
    .VS(VS),
    .CPU_HSYNC(HSYNC),
    .CPU_VSYNC(VSYNC),
    .CPU_FBLANK(FBLANK),
    .V(V),
    .RED(red),
    .GREEN(green),
    .BLUE(blue),

    .PALRAM_ADDR(PALRAM_ADDR),
    .PALRAM_DATA(PALRAM_DATA),

    .GAME(GAME),
    .FLIP(FLIP)
);

wire ym2151_cen, ym2151_cen2, oki_cen;
assign ym2151_cen = GAME == SNOWBRO2 ? CEN3p375 :
                    CEN3p375;
assign ym2151_cen2 = GAME == SNOWBRO2 ? CEN1p6875 :
                     CEN1p6875;
assign oki_cen = GAME == SNOWBRO2 ? CEN2p7 :
                 CEN2p7;

snowbro2_sound u_sound(
    .CLK(CLK),
    .CLK96(CLK96),
    .RESET(RESET),
    .RESET96(RESET96),
    .YM2151_CEN(ym2151_cen),
    .YM2151_CEN2(ym2151_cen2),
    .OKI_CEN(oki_cen),
    .PCM_CS(PCM_CS),
    .PCM_OK(PCM_OK),
    .PCM_ADDR(PCM_ADDR),
    .PCM_DOUT(PCM_DOUT),
    .left(snd_left),
    .right(snd_right),
    .sample(sample),
    .peak(peak),
    .YM2151_CS(YM2151_CS),
    .OKI_CS(OKI_CS),
    .YM2151_WE(YM2151_WE),
    .YM2151_WR_CMD(YM2151_WR_CMD),
    .OKI_WE(OKI_WE),
    .OKI_DIN(OKI_DIN),
    .YM2151_DIN(YM2151_DIN),
    .YM2151_DOUT(YM2151_DOUT),
    .OKI_DOUT(OKI_DOUT),
    .GAME(GAME),
    .FX_LEVEL(dip_fxlevel),
    .DIP_PAUSE(DIP_PAUSE),
    .OKI_BANK(OKI_BANK),
    .YM2151_INT(YM2151_INT)
);

//sdram
snowbro2_sdram u_sdram (
    .RESET(RESET96),
    .CLK(CLK96),
    .RESET48(RESET),
    .CLK48(CLK),
    .CLK_GFX(pxl_cen),

    //ROM loader
    .IOCTL_ADDR(ioctl_addr),
    .IOCTL_DOUT(ioctl_dout),
    .IOCTL_DIN(ioctl_din),
    .IOCTL_WR(ioctl_wr),
    .IOCTL_RAM(ioctl_ram),
    .PROG_ADDR(prog_addr),
    .PROG_DATA(prog_data),
    .PROG_MASK(prog_mask),
    .PROG_BA(prog_ba),
    .PROG_WE(prog_we),
    .PROG_RD(prog_rd),
    .PROG_RDY(prog_rdy),
    .DOWNLOADING(downloading),
    .DWNLD_BUSY(dwnld_busy),

    // Banks
    .BA0_ADDR(ba0_addr),
    .BA1_ADDR(ba1_addr),
    .BA2_ADDR(ba2_addr),
    .BA3_ADDR(ba3_addr),
    .BA_RD(ba_rd),
    .BA_WR(ba_wr),
    .BA0_DIN(ba0_din),
    .BA0_DIN_M(ba0_din_m),  // write mask
    .BA_ACK(ba_ack),
    .BA_DST(ba_dst),
    .BA_DOK(ba_dok),
    .BA_RDY(ba_rdy),
    .DATA_READ(data_read),

    //tiles
    .GFX_CS(GFX_CS),
    .GFX_OK(GFX_OK),
    .GFX0_ADDR(GFX0_ADDR),
    .GFX0_DOUT(GFX0_DOUT),

    .GFXSCR0_CS(GFXSCR0_CS),
    .GFXSCR0_OK(GFXSCR0_OK),
    .GFX0SCR0_ADDR(GFX0SCR0_ADDR),
    .GFX0SCR0_DOUT(GFX0SCR0_DOUT),

    .GFXSCR1_CS(GFXSCR1_CS),
    .GFXSCR1_OK(GFXSCR1_OK),
    .GFX0SCR1_ADDR(GFX0SCR1_ADDR),
    .GFX0SCR1_DOUT(GFX0SCR1_DOUT),

    .GFXSCR2_CS(GFXSCR2_CS),
    .GFXSCR2_OK(GFXSCR2_OK),
    .GFX0SCR2_ADDR(GFX0SCR2_ADDR),
    .GFX0SCR2_DOUT(GFX0SCR2_DOUT),

    //68k program
    .ROM68K_CS(ROM68K_CS),
    .ROM68K_OK(ROM68K_OK),
    .ROM68K_ADDR(ROM68K_ADDR),
    .ROM68K_DOUT(ROM68K_DOUT),

    //PCM data
    .PCM_CS(PCM_CS),
    .PCM_OK(PCM_OK),
    .PCM_ADDR(PCM_ADDR),
    .PCM_DOUT(PCM_DOUT),

    .GAME(GAME)
);

endmodule
